module state(
    input   wire   i_clk_sys,
    input   wire   i_rst_n,
    input   wire   i_
);
endmodule