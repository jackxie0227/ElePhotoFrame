module wifi(
    output CNT,
    output BOOT,
    output RESET
);

assign RESET = 1;
assign BOOT = 1;
assign CNT = 0;

endmodule
