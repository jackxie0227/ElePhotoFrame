/********************************************************************************
 * 模块名称: vga
 * 功能描述: VGA时序控制模块，生成800x600@60Hz的VGA时序信号
 *          产生水平同步信号(VGA_HS)、垂直同步信号(VGA_VS)和像素坐标
 * 
 * VGA 800x600@60Hz 时序参数:
 *   像素时钟频率: 40MHz
 *   水平扫描频率: 37.9KHz  
 *   垂直刷新频率: 60Hz
 *   
 * 水平时序: 1040个像素时钟周期
 *   同步脉冲: 120个时钟 | 后沿: 64个时钟 | 显示: 800个时钟 | 前沿: 56个时钟
 *   
 * 垂直时序: 660行
 *   同步脉冲: 6行 | 后沿: 23行 | 显示: 600行 | 前沿: 37行
 ********************************************************************************/
module vga(
    input  wire        clk,         // 像素时钟输入 (应为40MHz用于800x600@60Hz)
    output wire [9:0]  xpos,        // 当前像素X坐标 (0~799，有效显示区域)
    output wire [9:0]  ypos,        // 当前像素Y坐标 (0~599，有效显示区域)  
    output wire        VGA_HS,      // 水平同步信号 (负极性)
    output wire        VGA_VS       // 垂直同步信号 (负极性)
);

/************************VGA时序参数定义************************/
// 800x600@60Hz VGA标准时序参数
// 水平时序参数 (单位: 像素时钟周期)
/*************************************************************/
localparam H_TOTAL  = 1040;     // 水平总周期 = 120+64+800+56
localparam H_SYNC   = 120;      // 水平同步脉冲宽度
localparam H_BACK   = 64;       // 水平后沿时间  
localparam H_DISP   = 800;      // 水平显示时间
localparam H_FRONT  = 56;       // 水平前沿时间

/************************垂直时序参数定义************************/
// 垂直时序参数 (单位: 水平行数)
/*************************************************************/
localparam V_TOTAL  = 660;      // 垂直总周期 = 6+23+600+37  
localparam V_SYNC   = 6;        // 垂直同步脉冲宽度
localparam V_BACK   = 23;       // 垂直后沿时间
localparam V_DISP   = 600;      // 垂直显示时间
localparam V_FRONT  = 37;       // 垂直前沿时间

/************************显示区域边界计算************************/
// 用于确定有效显示区域的起始和结束位置
/*************************************************************/
localparam H_START  = H_SYNC + H_BACK;         // 水平显示区域起始位置 = 184
localparam H_END    = H_START + H_DISP;        // 水平显示区域结束位置 = 984
localparam V_START  = V_SYNC + V_BACK;         // 垂直显示区域起始位置 = 29  
localparam V_END    = V_START + V_DISP;        // 垂直显示区域结束位置 = 629

/************************扫描计数器************************/
// x_counter - 水平扫描计数器，范围0~1039
// y_counter - 垂直扫描计数器，范围0~659
/**********************************************************/
reg [11:0] x_counter;           // 水平扫描计数器 (12位，最大值1039)
reg [11:0] y_counter;           // 垂直扫描计数器 (12位，最大值659)

/************************计数器初始化************************/
// 系统上电时对扫描计数器进行初始化
// 避免仿真时出现未定义状态
/**********************************************************/
initial begin
    x_counter = 12'd0;
    y_counter = 12'd0;
end

/************************VGA扫描时序控制************************/
// posedge clk    在像素时钟的每个上升沿
// 
// 扫描顺序：
// 1. 水平扫描：从左到右逐像素扫描
// 2. 行扫描：完成一行后，转到下一行  
// 3. 场扫描：完成所有行后，从第一行重新开始
// 
// 计数器工作方式：
// - x_counter: 0→1→2→...→1039→0 (循环)
// - y_counter: 当x_counter=1039时递增，0→1→2→...→659→0
/*************************************************************/
always @(posedge clk) begin
    //****************水平扫描控制*****************/
    // 每个像素时钟周期递增水平计数器
    // 到达行末尾时清零并处理垂直计数
    /*******************************************/
    if (x_counter == H_TOTAL - 1) begin
        x_counter <= 12'd0;                 // 水平计数器清零，开始新行
        
        //****************垂直扫描控制*****************/
        // 每完成一行扫描递增垂直计数器
        // 到达帧末尾时清零，开始新帧
        /*******************************************/
        if (y_counter == V_TOTAL - 1) begin
            y_counter <= 12'd0;             // 垂直计数器清零，开始新帧
        end
        else begin
            y_counter <= y_counter + 1'b1;  // 垂直计数器递增，下一行
        end
    end
    else begin
        x_counter <= x_counter + 1'b1;      // 水平计数器递增，下一像素
    end
end

/************************VGA同步信号生成************************/
// VGA同步信号采用负极性
// VGA_HS: 水平同步信号，在同步脉冲期间为低电平
// VGA_VS: 垂直同步信号，在同步脉冲期间为低电平
// 
// 同步脉冲时序：
// - 水平同步: x_counter在0~119期间为低电平
// - 垂直同步: y_counter在0~5期间为低电平
/*************************************************************/
assign VGA_HS = ~(x_counter < H_SYNC);     // 水平同步信号（负极性）
assign VGA_VS = ~(y_counter < V_SYNC);     // 垂直同步信号（负极性）

/************************显示区域坐标输出************************/
// xpos, ypos: 当前像素在显示区域中的坐标
// 只在有效显示区域内输出有效坐标(0~799, 0~599)
// 在非显示区域坐标为负值，便于外部模块判断
// 
// 坐标计算:
// - xpos = x_counter - H_START  当x_counter∈[184,983]时，xpos∈[0,799]
// - ypos = y_counter - V_START  当y_counter∈[29,628]时，ypos∈[0,599]
/***************************************************************/
assign xpos = x_counter - H_START;         // X坐标偏移到显示区域
assign ypos = y_counter - V_START;         // Y坐标偏移到显示区域

/************************显示区域有效信号(可选)************************/
// 如果需要显示使能信号，可以取消以下注释
// 用于指示当前是否处于有效显示区域
/********************************************************************/
// wire display_valid;
// assign display_valid = (x_counter >= H_START && x_counter < H_END) &&
//                        (y_counter >= V_START && y_counter < V_END);

endmodule
