/********************************************************************************
 * 模块名称: clkdiv
 * 功能描述: 时钟分频模块，从50MHz输入时钟生成多个频率的输出时钟
 *          - clk_25m:  25MHz时钟，用于VGA显示或其他高频模块
 *          - clk_100k: 100KHz时钟，用于数码管扫描显示
 * 
 * 分频比计算:
 *   25MHz:  50MHz ÷ 2 = 25MHz   (计数范围: 0~1)
 *   100KHz: 50MHz ÷ 500 = 100KHz (计数范围: 0~249)
 ********************************************************************************/
module clkdiv(
    input  wire clk_50m,        // 输入50MHz系统时钟
    output reg  clk_25m,        // 输出25MHz时钟
    output reg  clk_100k        // 输出100KHz时钟
);

/************************时钟分频计数器************************/
// cnt_25m  - 25MHz时钟分频计数器，计数范围0~1
// cnt_100k - 100KHz时钟分频计数器，计数范围0~249  
/***********************************************************/
reg [0:0] cnt_25m;              // 25MHz分频计数器(1位)
reg [8:0] cnt_100k;             // 100KHz分频计数器(9位，最大值249)

/************************计数器初始化************************/
// 系统上电时对分频计数器进行初始化
// 避免仿真时出现未定义状态
/***********************************************************/
initial begin
    cnt_25m = 1'b0;
    cnt_100k = 9'd0;
    clk_25m = 1'b0;
    clk_100k = 1'b0;
end

/************************时钟分频逻辑************************/
// posedge clk_50m    在50MHz时钟的每个上升沿
// 
// 25MHz时钟生成：
// - 每2个50MHz时钟周期翻转一次输出
// - cnt_25m计数0~1，到1时翻转clk_25m并清零计数器
// 
// 100KHz时钟生成：
// - 每250个50MHz时钟周期翻转一次输出  
// - cnt_100k计数0~249，到249时翻转clk_100k并清零计数器
/***********************************************************/
always @(posedge clk_50m) begin
    //****************25MHz时钟生成*****************/
    // 分频比：50MHz ÷ 2 = 25MHz
    // 计数周期：每2个时钟周期翻转一次输出
    // 占空比：50% (高电平1个周期，低电平1个周期)
    /*********************************************/
    if (cnt_25m == 1'b1) begin
        clk_25m <= ~clk_25m;        // 翻转25MHz时钟输出
        cnt_25m <= 1'b0;            // 计数器清零重新开始
    end
    else begin
        cnt_25m <= cnt_25m + 1'b1;  // 计数器递增
    end
    
    //****************100KHz时钟生成*****************/
    // 分频比：50MHz ÷ 500 = 100KHz  
    // 计数周期：每250个时钟周期翻转一次输出
    // 占空比：50% (高电平250个周期，低电平250个周期)
    /***********************************************/
    if (cnt_100k == 9'd249) begin
        clk_100k <= ~clk_100k;      // 翻转100KHz时钟输出
        cnt_100k <= 9'd0;           // 计数器清零重新开始
    end
    else begin
        cnt_100k <= cnt_100k + 1'b1; // 计数器递增
    end
end

endmodule
