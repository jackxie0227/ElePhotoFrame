/********************************************************************************
 * 模块名称: clkdiv
 * 功能描述: 时钟分频模块，从50MHz输入时钟生成多个频率的输出时钟
 *          - clk_5m:   5MHz时钟，用于特定模块
 *          - clk_100k: 100KHz时钟，用于数码管扫描显示
 * 
 * 分频比计算:
 *   5MHz:   50MHz ÷ 10 = 5MHz   (计数范围: 0~4)
 *   100KHz: 50MHz ÷ 500 = 100KHz (计数范围: 0~249)
 ********************************************************************************/
module clkdiv(
    input  wire clk_50m,        // 输入50MHz系统时钟
    output reg  clk_5m,         // 输出5MHz时钟
    output reg  clk_100k        // 输出100KHz时钟
);

/************************时钟分频计数器************************/
// cnt_5m   - 5MHz时钟分频计数器，计数范围0~4
// cnt_100k - 100KHz时钟分频计数器，计数范围0~249  
/***********************************************************/
reg [2:0] cnt_5m;               // 5MHz分频计数器(3位)
reg [8:0] cnt_100k;             // 100KHz分频计数器(9位，最大值249)

/************************计数器初始化************************/
// 系统上电时对分频计数器进行初始化
// 避免仿真时出现未定义状态
/***********************************************************/
initial begin
    cnt_5m = 3'd0;
    cnt_100k = 9'd0;
    clk_5m = 1'b0;
    clk_100k = 1'b0;
end

/************************时钟分频逻辑************************/
// posedge clk_50m    在50MHz时钟的每个上升沿
// 
// 5MHz时钟生成：
// - 每10个50MHz时钟周期翻转一次输出
// - cnt_5m计数0~4，到4时翻转clk_5m并清零计数器
// 
// 100KHz时钟生成：
// - 每250个50MHz时钟周期翻转一次输出  
// - cnt_100k计数0~249，到249时翻转clk_100k并清零计数器
/***********************************************************/
always @(posedge clk_50m) begin
    //****************5MHz时钟生成*****************/
    // 分频比：50MHz ÷ 10 = 5MHz
    // 计数周期：每5个时钟周期翻转一次输出
    // 占空比：50% (高电平5个周期，低电平5个周期)
    /*********************************************/
    if (cnt_5m == 3'd4) begin
        clk_5m <= ~clk_5m;          // 翻转5MHz时钟输出
        cnt_5m <= 3'd0;             // 计数器清零重新开始
    end
    else begin
        cnt_5m <= cnt_5m + 3'd1;    // 计数器递增
    end
    
    //****************100KHz时钟生成*****************/
    // 分频比：50MHz ÷ 500 = 100KHz  
    // 计数周期：每250个时钟周期翻转一次输出
    // 占空比：50% (高电平250个周期，低电平250个周期)
    /***********************************************/
    if (cnt_100k == 9'd249) begin
        clk_100k <= ~clk_100k;      // 翻转100KHz时钟输出
        cnt_100k <= 9'd0;           // 计数器清零重新开始
    end
    else begin
        cnt_100k <= cnt_100k + 1'b1; // 计数器递增
    end
end

endmodule
